LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MYFIFO_1 IS
	PORT ( DATAIN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		EN,CLK,RST : IN STD_LOGIC ;
		W : IN STD_LOGIC;
		DATAOUT : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0);
		RED : OUT STD_LOGIC);
END MYFIFO_1;

ARCHITECTURE BEHAVIORAL OF MYFIFO_1 IS

SIGNAL WPTR, RPTR : STD_LOGIC_VECTOR(3 DOWNTO 0);
TYPE FIFO IS ARRAY(15 DOWNTO 00) OF STD_LOGIC_VECTOR(07 DOWNTO 00);
SIGNAL MEM:FIFO;

BEGIN

PROCESS(CLK,RST)
BEGIN
	IF RST = '1' THEN
		WPTR <= "0000" ;
		RPTR <= "0000" ;
		RED <= '0' ;
	ELSE IF(CLK' EVENT AND CLK='1') THEN
		IF(EN = '1') THEN
			IF(W = '1') THEN               -- Write Operation
				IF(WPTR < "1111") THEN
				 	MEM(CONV_INTEGER(WPTR)) <= DATAIN;
					WPTR <= WPTR + 1 ;
				ELSE
					RED <= '1' ;   -- Memory Full Warning
				END IF ;
			ELSE                           -- Read Operation
				IF(RPTR < WPTR) THEN
					RED <= '0';
					DATAOUT <= MEM(CONV_INTEGER(RPTR));
					RPTR <= RPTR + 1;
				ELSE
					RED <= '1' ;   -- Empty Memory Warning
					DATAOUT <= "00000000" ;
				END IF ;
			END IF ;
		END iF ;
	END IF ;
END IF ;
END PROCESS ;
END BEHAVIORAL ;




 
		
